Biolek R2 Model for a Bipolar Threshold Memristive Device
********************************************************************************
* Connections:
* p - top electrode
* n - bottom electrode
* x - External connection to plot state variable that is not used otherwise
********************************************************************************
.SUBCKT BiolekR2 p n PARAMS: xinit=0.11
********************************************************************************
* Device Constants
*********************************************************************************
.PARAMS Ron=1k Roff=10k Rinit=(Ron+Roff)/2 Beta=1e13 Vt=4.6V b1=10u b2=10u x0={xinit}

.PARAM Cval=1
********************************************************************************
* Theta Function
********************************************************************************
.FUNC theta(x, b)  {1 / (1 + EXP(-x / b))}
********************************************************************************
* Gamma Function
********************************************************************************
.FUNC gamma(x, b)  {x * ({theta(x, b)} - {theta(-x, b)})}
