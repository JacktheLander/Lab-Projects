Dual RC ladder
********************************************************************************
R1 int in 10k
V1 in 0 dc 0 ac 1
R2 out int 1k
C1 int 0 1u
C2 out 0 100n
.ac dec 10 1 100k
.control
run
.endc
.end
